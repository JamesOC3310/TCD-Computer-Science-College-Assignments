----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12/20/2021 04:32:14 PM
-- Design Name: 
-- Module Name: ControlMemory_20332090 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--use IEEE.STD_LOGIC_ARITH.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ControlMemory_20332090 is
  Port ( IN_CAR : in std_logic_vector(16 downto 0);
         FL : out std_logic; -- 0
         RZ : out std_logic; -- 1
         RN : out std_logic; -- 2
         RC : out std_logic; -- 3
         RV : out std_logic; -- 4
         MW : out std_logic; -- 5
         MM : out std_logic; -- 6
         RW : out std_logic; -- 7
         MD : out std_logic; -- 8
         FS : out std_logic_vector(4 downto 0); -- 9 to 13
         MB : out std_logic; -- 14
         TB : out std_logic; -- 15
         TA : out std_logic; -- 16
         TD : out std_logic; -- 17
         PL : out std_logic; -- 18
         PI : out std_logic; -- 19
         IL : out std_logic; -- 20
         MC : out std_logic; -- 21
         MS : out std_logic_vector(2 downto 0); -- 22 to 24
         NA : out std_logic_vector(16 downto 0) -- 25 to 41
 );
end ControlMemory_20332090;

architecture Behavioral of ControlMemory_20332090 is

        -- we will use the least significant 8 bit of the IN_CAR - array(0 to 255)
        type mem_array is array(0 to 255) of std_logic_vector(41 downto 0);
        
   -- initialise the control memory
        signal control_mem : mem_array := (
        -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address | MS | M| I| P| P| T| T| T| M| FS |M|R|M|M|R|R|R|R|F|vioral;
        -- | Next Address | MS | C| L| I| L| D| A| B| B| FS |D|W|M|W|V|C|N|Z|L|
        -- "00000000000000000 000 0 0 0 0 0 0 0 0 00000 0 0 0 0 0 0 0 0 0"
       "000000000000000000000000000000000000000000",-- 00
       "000000000000000000000000000000000000000000",-- 01 XOR R[DR] <- R[SA] XOR R[SB]
       --"000000000001001111110000100000000010000000",-- 02 LD  R[DR] <- M[R[SA]]
       --"000000000110000000010000000011000010000000",-- 03 srn R[DR] <- n R[SA] sr R[SB]
       --"000000000110000000010000000000000110000000",-- 04 INC R[DR] <- R[SA] + 1
       --"000000000000001010000000000000000000000000",-- 05
       --"000000000000001100000000000000000000000000",-- 06
       --"000000000000001110000000000000000000000000",-- 07
       ---- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
       ---- | Next Address | MS | M| I| P| P| T| T| T| M| FS |M|R|M|M|R|R|R|R|F|
       ---- | Next Address | MS | C| L| I| L| D| A| B| B| FS |D|W|M|W|V|C|N|Z|L|
       ---- "00000000000000000 000 0 0 0 0 0 0 0 0 00000 0 0 0 0 0 0 0 0 0"
       --"000000000000010000000000000000000000000000",-- 08
       --"000000000000010010000000000000000000000000",-- 09
       --"000000000000010100000000000000000000000000",-- 0A
       --"000000000000010110000000000000000000000000",-- 0B
       --"000000000000011000000000000000000000000000",-- 0C
       --"000000000000011010000000000000000000000000",-- 0D
       --"000000000000011100000000000000000000000000",-- 0E
       --"000000000000011110000000000000000000000000",-- 0F
       ---- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
       ---- | Next Address | MS | M| I| P| P| T| T| T| M| FS |M|R|M|M|R|R|R|R|F|
       ---- | Next Address | MS | C| L| I| L| D| A| B| B| FS |D|W|M|W|V|C|N|Z|L|
       ---- "00000000000000000 000 0 0 0 0 0 0 0 0 00000 0 0 0 0 0 0 0 0 0"
       --"000000000000100000000000000000000000000000",-- 10
       --"000000000000100010000000000000000000000000",-- 11
       --"000000000000100100000000000000000000000000",-- 12
       --"000000000000100110000000000000000000000000",-- 13
       --"000000000000101000000000000000000000000000",-- 14
       --"000000000000101010000000000000000000000000",-- 15
       --"000000000000101100000000000000000000000000",-- 16
       --"000000000000101110000000000000000000000000",-- 17
       --
       --"000000000000110000000000000000000000000000",
       --"000000000000110010000000000000000000000000",
       --"000000000000110100000000000000000000000000",
       --"000000000000110110000000000000000000000000",
       
        
      
        -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address | MS | M| I| P| P| T| T| T| M| FS |M|R|M|M|R|R|R|R|F|
        -- | Next Address | MS | C| L| I| L| D| A| B| B| FS |D|W|M|W|V|C|N|Z|L|
        -- "00000000000000000 000 0 0 0 0 0 0 0 0 00000 0 0 0 0 0 0 0 0 0"
      --  "000000000111110000000000000000000000000000",-- F8
      --"000000000111110010000000000000000000000000",-- F9
      --"000000000111110100000000000000000000000000",-- FA
      --"000000000111110110000000000000000000000000",-- FB
      --"000000000111111000000000000000000000000000",-- FC
      --"000000000111111010000000000000000000000000",-- FD
      --"000000000111111100000000000000000000000000",-- FE
      --"000000000111111110000000000000000000000000" -- FF
      
     "000000000010110100000000000000000000000000",
     "000000000101101100000000000000000000000000",
     "000000000101110000000000000000000000000000",
     "000000000101110100000000000000000000000000",
     "000000000101111000000000000000000000000000",
     "000000000101111100000000000000000000000000",
     "000000000110000000000000000000000000000000",
     "000000000110000100000000000000000000000000",
     "000000000110001000000000000000000000000000",
     "000000000110001100000000000000000000000000",
     "000000000110010000000000000000000000000000",
     "000000000110010100000000000000000000000000",
     "000000000110011000000000000000000000000000",
     "000000000110011100000000000000000000000000",
     "000000000110100000000000000000000000000000",
     "000000000110100100000000000000000000000000",
     "000000000110101000000000000000000000000000",
     "000000000110101100000000000000000000000000",
     "000000000110110000000000000000000000000000",
     "000000000110110100000000000000000000000000",
     "000000000110111000000000000000000000000000",
     "000000000110111100000000000000000000000000",
     "000000000111000000000000000000000000000000",
     "000000000111000100000000000000000000000000",
     "000000000111001000000000000000000000000000",
     "000000000111001100000000000000000000000000",
     "000000000111010000000000000000000000000000",
     "000000000111010100000000000000000000000000",
     "000000000111011000000000000000000000000000",
     "000000000111011100000000000000000000000000",
     "000000000111100000000000000000000000000000",
     "000000000111100100000000000000000000000000",
     "000000000111101000000000000000000000000000",
     "000000000111101100000000000000000000000000",
     "000000000111110000000000000000000000000000",
     "000000000111110100000000000000000000000000",
     "000000000111111000000000000000000000000000",
     "000000000111111100000000000000000000000000",
     "000000001000000000000000000000000000000000",
     "000000001000000100000000000000000000000000",
     "000000001000001000000000000000000000000000",
     "000000001000001100000000000000000000000000",
     "000000001000010000000000000000000000000000",
     "000000001000010100000000000000000000000000",
     "000000001000011000000000000000000000000000",
     "000000001000011100000000000000000000000000",
     "000000001000100000000000000000000000000000",
     "000000001000100100000000000000000000000000",
     "000000001000101000000000000000000000000000",
     "000000001000101100000000000000000000000000",
     "000000001000110000000000000000000000000000",
     "000000001000110100000000000000000000000000",
     "000000001000111000000000000000000000000000",
     "000000001000111100000000000000000000000000",
     "000000001001000000000000000000000000000000",
     "000000001001000100000000000000000000000000",
     "000000001001001000000000000000000000000000",
     "000000001001001100000000000000000000000000",
     "000000001001010000000000000000000000000000",
     "000000001001010100000000000000000000000000",
     "000000001001011000000000000000000000000000",
     "000000001001011100000000000000000000000000",
     "000000001001100000000000000000000000000000",
     "000000001001100100000000000000000000000000",
     "000000001001101000000000000000000000000000",
     "000000001001101100000000000000000000000000",
     "000000001001110000000000000000000000000000",
     "000000001001110100000000000000000000000000",
     "000000001001111000000000000000000000000000",
     "000000001001111100000000000000000000000000",
     "000000001010000000000000000000000000000000",
     "000000001010000100000000000000000000000000",
     "000000001010001000000000000000000000000000",
     "000000001010001100000000000000000000000000",
     "000000001010010000000000000000000000000000",
     "000000001010010100000000000000000000000000",
     "000000001010011000000000000000000000000000",
     "000000001010011100000000000000000000000000",
     "000000001010100000000000000000000000000000",
     "000000001010100100000000000000000000000000",
     "000000001010101000000000000000000000000000",
     "000000001010101100000000000000000000000000",
     "000000001010110000000000000000000000000000",
     "000000001010110100000000000000000000000000",
     "000000001010111000000000000000000000000000",
     "000000001010111100000000000000000000000000",
     "000000001011000000000000000000000000000000",
     "000000001011000100000000000000000000000000",
     "000000001011001000000000000000000000000000",
     "000000001011001100000000000000000000000000",
     "000000001011010000000000000000000000000000",
     "000000001011010100000000000000000000000000",
     "000000001011011000000000000000000000000000",
     "000000001011011100000000000000000000000000",
     "000000001011100000000000000000000000000000",
     "000000001011100100000000000000000000000000",
     "000000001011101000000000000000000000000000",
     "000000001011101100000000000000000000000000",
     "000000001011110000000000000000000000000000",
     "000000001011110100000000000000000000000000",
     "000000001011111000000000000000000000000000",
     "000000001011111100000000000000000000000000",
     "000000001100000000000000000000000000000000",
     "000000001100000100000000000000000000000000",
     "000000001100001000000000000000000000000000",
     "000000001100001100000000000000000000000000",
     "000000001100010000000000000000000000000000",
     "000000001100010100000000000000000000000000",
     "000000001100011000000000000000000000000000",
     "000000001100011100000000000000000000000000",
     "000000001100100000000000000000000000000000",
     "000000001100100100000000000000000000000000",
     "000000001100101000000000000000000000000000",
     "000000001100101100000000000000000000000000",
     "000000001100110000000000000000000000000000",
     "000000001100110100000000000000000000000000",
     "000000001100111000000000000000000000000000",
     "000000001100111100000000000000000000000000",
     "000000001101000000000000000000000000000000",
     "000000001101000100000000000000000000000000",
     "000000001101001000000000000000000000000000",
     "000000001101001100000000000000000000000000",
     "000000001101010000000000000000000000000000",
     "000000001101010100000000000000000000000000",
     "000000001101011000000000000000000000000000",
     "000000001101011100000000000000000000000000",
     "000000001101100000000000000000000000000000",
     "000000001101100100000000000000000000000000",
     "000000001101101000000000000000000000000000",
     "000000001101101100000000000000000000000000",
     "000000001101110000000000000000000000000000",
     "000000001101110100000000000000000000000000",
     "000000001101111000000000000000000000000000",
     "000000001101111100000000000000000000000000",
     "000000001110000000000000000000000000000000",
     "000000001110000100000000000000000000000000",
     "000000001110001000000000000000000000000000",
     "000000001110001100000000000000000000000000",
     "000000001110010000000000000000000000000000",
     "000000001110010100000000000000000000000000",
     "000000001110011000000000000000000000000000",
     "000000001110011100000000000000000000000000",
     "000000001110100000000000000000000000000000",
     "000000001110100100000000000000000000000000",
     "000000001110101000000000000000000000000000",
     "000000001110101100000000000000000000000000",
     "000000001110110000000000000000000000000000",
     "000000001110110100000000000000000000000000",
     "000000001110111000000000000000000000000000",
     "000000001110111100000000000000000000000000",
     "000000001111000000000000000000000000000000",
     "000000001111000100000000000000000000000000",
     "000000001111001000000000000000000000000000",
     "000000001111001100000000000000000000000000",
     "000000001111010000000000000000000000000000",
     "000000001111010100000000000000000000000000",
     "000000001111011000000000000000000000000000",
     "000000001111011100000000000000000000000000",
     "000000001111100000000000000000000000000000",
     "000000001111100100000000000000000000000000",
     "000000001111101000000000000000000000000000",
     "000000001111101100000000000000000000000000",
     "000000001111110000000000000000000000000000",
     "000000001111110100000000000000000000000000",
     "000000001111111000000000000000000000000000",
     "000000001111111100000000000000000000000000",
     "000000010000000000000000000000000000000000",
     "000000010000000100000000000000000000000000",
     "000000010000001000000000000000000000000000",
     "000000010000001100000000000000000000000000",
     "000000010000010000000000000000000000000000",
     "000000010000010100000000000000000000000000",
     "000000010000011000000000000000000000000000",
     "000000010000011100000000000000000000000000",
     "000000010000100000000000000000000000000000",
     "000000010000100100000000000000000000000000",
     "000000010000101000000000000000000000000000",
     "000000010000101100000000000000000000000000",
     "000000010000110000000000000000000000000000",
     "000000010000110100000000000000000000000000",
     "000000010000111000000000000000000000000000",
     "000000010000111100000000000000000000000000",
     "000000010001000000000000000000000000000000",
     "000000010001000100000000000000000000000000",
     "000000010001001000000000000000000000000000",
     "000000010001001100000000000000000000000000",
     "000000010001010000000000000000000000000000",
     "000000010001010100000000000000000000000000",
     "000000010001011000000000000000000000000000",
     "000000010001011100000000000000000000000000",
     "000000010001100000000000000000000000000000",
     "000000010001100100000000000000000000000000",
     "000000010001101000000000000000000000000000",
     "000000010001101100000000000000000000000000",
     "000000010001110000000000000000000000000000",
     "000000010001110100000000000000000000000000",
     "000000010001111000000000000000000000000000",
     "000000010001111100000000000000000000000000",
     "000000010010000000000000000000000000000000",
     "000000010010000100000000000000000000000000",
     "000000010010001000000000000000000000000000",
     "000000010010001100000000000000000000000000",
     "000000010010010000000000000000000000000000",
     "000000010010010100000000000000000000000000",
     "000000010010011000000000000000000000000000",
     "000000010010011100000000000000000000000000",
     "000000010010100000000000000000000000000000",
     "000000010010100100000000000000000000000000",
     "000000010010101000000000000000000000000000",
     "000000010010101100000000000000000000000000",
     "000000010010110000000000000000000000000000",
     "000000010010110100000000000000000000000000",
     "000000010010111000000000000000000000000000",
     "000000010010111100000000000000000000000000",
     "000000010011000000000000000000000000000000",
     "000000010011000100000000000000000000000000",
     "000000010011001000000000000000000000000000",
     "000000010011001100000000000000000000000000",
     "000000010011010000000000000000000000000000",
     "000000010011010100000000000000000000000000",
     "000000010011011000000000000000000000000000",
     "000000010011011100000000000000000000000000",
     "000000010011100000000000000000000000000000",
     "000000010011100100000000000000000000000000",
     "000000010011101000000000000000000000000000",
     "000000010011101100000000000000000000000000",
     "000000010011110000000000000000000000000000",
     "000000010011110100000000000000000000000000",
     "000000010011111000000000000000000000000000",
     "000000010011111100000000000000000000000000",
     "000000010100000000000000000000000000000000",
     "000000010100000100000000000000000000000000",
     "000000010100001000000000000000000000000000",
     "000000010100001100000000000000000000000000",
     "000000010100010000000000000000000000000000",
     "000000010100010100000000000000000000000000",
     "000000010100011000000000000000000000000000",
     "000000010100011100000000000000000000000000",
     "000000010100100000000000000000000000000000",
     "000000010100100100000000000000000000000000",
     "000000010100101000000000000000000000000000",
     "000000010100101100000000000000000000000000",
     "000000010100110000000000000000000000000000",
     "000000010100110100000000000000000000000000",
     "000000010100111000000000000000000000000000",
     "000000010100111100000000000000000000000000",
     "000000010101000000000000000000000000000000",
     "000000010101000100000000000000000000000000",
     "000000010101001000000000000000000000000000",
     "000000010101001100000000000000000000000000",
     "000000010101010000000000000000000000000000",
     "000000010101010100000000000000000000000000",
     "000000010101011000000000000000000000000000",
     "000000010101011100000000000000000000000000"
     --"000000010101100000000000000000000000000000",
     --"000000010101100100000000000000000000000000"    
       );
        
        signal content_at_address : std_logic_vector(41 downto 0); 
begin
        content_at_address <= control_mem(to_integer(unsigned(IN_CAR(8 downto 0)))) after 2ns;
        FL <= content_at_address(0); -- 0
        RZ <= content_at_address(1); -- 1
        RN <= content_at_address(2); -- 2
        RC <= content_at_address(3); -- 3
        RV <= content_at_address(4); -- 4
        MW <= content_at_address(5); -- 5
        MM <= content_at_address(6); -- 6
        RW <= content_at_address(7); -- 7
        MD <= content_at_address(8); -- 8
        FS <= content_at_address(13 downto 9); -- 9 to 13
        MB <= content_at_address(14); -- 14
        
        TB <= content_at_address(15); -- 15
        TA <= content_at_address(16); -- 16
        TD <= content_at_address(17); -- 17
        PL <= content_at_address(18); -- 18
        PI <= content_at_address(19); -- 19
        IL <= content_at_address(20); -- 20
        MC <= content_at_address(21); -- 21
        MS <= content_at_address(24 downto 22); -- 22 to 24
        NA <= content_at_address(41 downto 25); -- 25 to 41
        

end Behavioral;